../../test_cases/ispd19/ispd19_test1/ispd19_test1.input.lef